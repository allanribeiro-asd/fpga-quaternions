library verilog;
use verilog.vl_types.all;
entity system_0_rsp_xbar_mux_001 is
    port(
        sink0_valid     : in     vl_logic;
        sink0_data      : in     vl_logic_vector(101 downto 0);
        sink0_channel   : in     vl_logic_vector(23 downto 0);
        sink0_startofpacket: in     vl_logic;
        sink0_endofpacket: in     vl_logic;
        sink0_ready     : out    vl_logic;
        sink1_valid     : in     vl_logic;
        sink1_data      : in     vl_logic_vector(101 downto 0);
        sink1_channel   : in     vl_logic_vector(23 downto 0);
        sink1_startofpacket: in     vl_logic;
        sink1_endofpacket: in     vl_logic;
        sink1_ready     : out    vl_logic;
        sink2_valid     : in     vl_logic;
        sink2_data      : in     vl_logic_vector(101 downto 0);
        sink2_channel   : in     vl_logic_vector(23 downto 0);
        sink2_startofpacket: in     vl_logic;
        sink2_endofpacket: in     vl_logic;
        sink2_ready     : out    vl_logic;
        sink3_valid     : in     vl_logic;
        sink3_data      : in     vl_logic_vector(101 downto 0);
        sink3_channel   : in     vl_logic_vector(23 downto 0);
        sink3_startofpacket: in     vl_logic;
        sink3_endofpacket: in     vl_logic;
        sink3_ready     : out    vl_logic;
        sink4_valid     : in     vl_logic;
        sink4_data      : in     vl_logic_vector(101 downto 0);
        sink4_channel   : in     vl_logic_vector(23 downto 0);
        sink4_startofpacket: in     vl_logic;
        sink4_endofpacket: in     vl_logic;
        sink4_ready     : out    vl_logic;
        sink5_valid     : in     vl_logic;
        sink5_data      : in     vl_logic_vector(101 downto 0);
        sink5_channel   : in     vl_logic_vector(23 downto 0);
        sink5_startofpacket: in     vl_logic;
        sink5_endofpacket: in     vl_logic;
        sink5_ready     : out    vl_logic;
        sink6_valid     : in     vl_logic;
        sink6_data      : in     vl_logic_vector(101 downto 0);
        sink6_channel   : in     vl_logic_vector(23 downto 0);
        sink6_startofpacket: in     vl_logic;
        sink6_endofpacket: in     vl_logic;
        sink6_ready     : out    vl_logic;
        sink7_valid     : in     vl_logic;
        sink7_data      : in     vl_logic_vector(101 downto 0);
        sink7_channel   : in     vl_logic_vector(23 downto 0);
        sink7_startofpacket: in     vl_logic;
        sink7_endofpacket: in     vl_logic;
        sink7_ready     : out    vl_logic;
        sink8_valid     : in     vl_logic;
        sink8_data      : in     vl_logic_vector(101 downto 0);
        sink8_channel   : in     vl_logic_vector(23 downto 0);
        sink8_startofpacket: in     vl_logic;
        sink8_endofpacket: in     vl_logic;
        sink8_ready     : out    vl_logic;
        sink9_valid     : in     vl_logic;
        sink9_data      : in     vl_logic_vector(101 downto 0);
        sink9_channel   : in     vl_logic_vector(23 downto 0);
        sink9_startofpacket: in     vl_logic;
        sink9_endofpacket: in     vl_logic;
        sink9_ready     : out    vl_logic;
        sink10_valid    : in     vl_logic;
        sink10_data     : in     vl_logic_vector(101 downto 0);
        sink10_channel  : in     vl_logic_vector(23 downto 0);
        sink10_startofpacket: in     vl_logic;
        sink10_endofpacket: in     vl_logic;
        sink10_ready    : out    vl_logic;
        sink11_valid    : in     vl_logic;
        sink11_data     : in     vl_logic_vector(101 downto 0);
        sink11_channel  : in     vl_logic_vector(23 downto 0);
        sink11_startofpacket: in     vl_logic;
        sink11_endofpacket: in     vl_logic;
        sink11_ready    : out    vl_logic;
        sink12_valid    : in     vl_logic;
        sink12_data     : in     vl_logic_vector(101 downto 0);
        sink12_channel  : in     vl_logic_vector(23 downto 0);
        sink12_startofpacket: in     vl_logic;
        sink12_endofpacket: in     vl_logic;
        sink12_ready    : out    vl_logic;
        sink13_valid    : in     vl_logic;
        sink13_data     : in     vl_logic_vector(101 downto 0);
        sink13_channel  : in     vl_logic_vector(23 downto 0);
        sink13_startofpacket: in     vl_logic;
        sink13_endofpacket: in     vl_logic;
        sink13_ready    : out    vl_logic;
        sink14_valid    : in     vl_logic;
        sink14_data     : in     vl_logic_vector(101 downto 0);
        sink14_channel  : in     vl_logic_vector(23 downto 0);
        sink14_startofpacket: in     vl_logic;
        sink14_endofpacket: in     vl_logic;
        sink14_ready    : out    vl_logic;
        sink15_valid    : in     vl_logic;
        sink15_data     : in     vl_logic_vector(101 downto 0);
        sink15_channel  : in     vl_logic_vector(23 downto 0);
        sink15_startofpacket: in     vl_logic;
        sink15_endofpacket: in     vl_logic;
        sink15_ready    : out    vl_logic;
        sink16_valid    : in     vl_logic;
        sink16_data     : in     vl_logic_vector(101 downto 0);
        sink16_channel  : in     vl_logic_vector(23 downto 0);
        sink16_startofpacket: in     vl_logic;
        sink16_endofpacket: in     vl_logic;
        sink16_ready    : out    vl_logic;
        sink17_valid    : in     vl_logic;
        sink17_data     : in     vl_logic_vector(101 downto 0);
        sink17_channel  : in     vl_logic_vector(23 downto 0);
        sink17_startofpacket: in     vl_logic;
        sink17_endofpacket: in     vl_logic;
        sink17_ready    : out    vl_logic;
        sink18_valid    : in     vl_logic;
        sink18_data     : in     vl_logic_vector(101 downto 0);
        sink18_channel  : in     vl_logic_vector(23 downto 0);
        sink18_startofpacket: in     vl_logic;
        sink18_endofpacket: in     vl_logic;
        sink18_ready    : out    vl_logic;
        sink19_valid    : in     vl_logic;
        sink19_data     : in     vl_logic_vector(101 downto 0);
        sink19_channel  : in     vl_logic_vector(23 downto 0);
        sink19_startofpacket: in     vl_logic;
        sink19_endofpacket: in     vl_logic;
        sink19_ready    : out    vl_logic;
        sink20_valid    : in     vl_logic;
        sink20_data     : in     vl_logic_vector(101 downto 0);
        sink20_channel  : in     vl_logic_vector(23 downto 0);
        sink20_startofpacket: in     vl_logic;
        sink20_endofpacket: in     vl_logic;
        sink20_ready    : out    vl_logic;
        sink21_valid    : in     vl_logic;
        sink21_data     : in     vl_logic_vector(101 downto 0);
        sink21_channel  : in     vl_logic_vector(23 downto 0);
        sink21_startofpacket: in     vl_logic;
        sink21_endofpacket: in     vl_logic;
        sink21_ready    : out    vl_logic;
        sink22_valid    : in     vl_logic;
        sink22_data     : in     vl_logic_vector(101 downto 0);
        sink22_channel  : in     vl_logic_vector(23 downto 0);
        sink22_startofpacket: in     vl_logic;
        sink22_endofpacket: in     vl_logic;
        sink22_ready    : out    vl_logic;
        sink23_valid    : in     vl_logic;
        sink23_data     : in     vl_logic_vector(101 downto 0);
        sink23_channel  : in     vl_logic_vector(23 downto 0);
        sink23_startofpacket: in     vl_logic;
        sink23_endofpacket: in     vl_logic;
        sink23_ready    : out    vl_logic;
        src_valid       : out    vl_logic;
        src_data        : out    vl_logic_vector(101 downto 0);
        src_channel     : out    vl_logic_vector(23 downto 0);
        src_startofpacket: out    vl_logic;
        src_endofpacket : out    vl_logic;
        src_ready       : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end system_0_rsp_xbar_mux_001;
