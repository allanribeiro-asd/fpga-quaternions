library verilog;
use verilog.vl_types.all;
entity system_0_cfi_flash_0 is
    generic(
        TCM_ADDRESS_W   : integer := 22;
        TCM_DATA_W      : integer := 8;
        TCM_BYTEENABLE_W: integer := 1;
        TCM_READ_WAIT   : integer := 160;
        TCM_WRITE_WAIT  : integer := 160;
        TCM_SETUP_WAIT  : integer := 40;
        TCM_DATA_HOLD   : integer := 40;
        TCM_TURNAROUND_TIME: integer := 2;
        TCM_TIMING_UNITS: integer := 0;
        TCM_READLATENCY : integer := 2;
        TCM_SYMBOLS_PER_WORD: integer := 1;
        USE_READDATA    : integer := 1;
        USE_WRITEDATA   : integer := 1;
        USE_READ        : integer := 1;
        USE_WRITE       : integer := 1;
        USE_BYTEENABLE  : integer := 0;
        USE_CHIPSELECT  : integer := 1;
        USE_LOCK        : integer := 0;
        USE_ADDRESS     : integer := 1;
        USE_WAITREQUEST : integer := 0;
        USE_WRITEBYTEENABLE: integer := 0;
        USE_OUTPUTENABLE: integer := 0;
        USE_RESETREQUEST: integer := 0;
        USE_IRQ         : integer := 0;
        USE_RESET_OUTPUT: integer := 0;
        ACTIVE_LOW_READ : integer := 1;
        ACTIVE_LOW_LOCK : integer := 0;
        ACTIVE_LOW_WRITE: integer := 1;
        ACTIVE_LOW_CHIPSELECT: integer := 1;
        ACTIVE_LOW_BYTEENABLE: integer := 0;
        ACTIVE_LOW_OUTPUTENABLE: integer := 0;
        ACTIVE_LOW_WRITEBYTEENABLE: integer := 0;
        ACTIVE_LOW_WAITREQUEST: integer := 0;
        ACTIVE_LOW_BEGINTRANSFER: integer := 0;
        CHIPSELECT_THROUGH_READLATENCY: integer := 0
    );
    port(
        clk_clk         : in     vl_logic;
        reset_reset     : in     vl_logic;
        uas_address     : in     vl_logic_vector(21 downto 0);
        uas_burstcount  : in     vl_logic_vector(0 downto 0);
        uas_read        : in     vl_logic;
        uas_write       : in     vl_logic;
        uas_waitrequest : out    vl_logic;
        uas_readdatavalid: out    vl_logic;
        uas_byteenable  : in     vl_logic_vector(0 downto 0);
        uas_readdata    : out    vl_logic_vector(7 downto 0);
        uas_writedata   : in     vl_logic_vector(7 downto 0);
        uas_lock        : in     vl_logic;
        uas_debugaccess : in     vl_logic;
        tcm_write_n_out : out    vl_logic;
        tcm_read_n_out  : out    vl_logic;
        tcm_chipselect_n_out: out    vl_logic;
        tcm_request     : out    vl_logic;
        tcm_grant       : in     vl_logic;
        tcm_address_out : out    vl_logic_vector(21 downto 0);
        tcm_data_out    : out    vl_logic_vector(7 downto 0);
        tcm_data_outen  : out    vl_logic;
        tcm_data_in     : in     vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TCM_ADDRESS_W : constant is 1;
    attribute mti_svvh_generic_type of TCM_DATA_W : constant is 1;
    attribute mti_svvh_generic_type of TCM_BYTEENABLE_W : constant is 1;
    attribute mti_svvh_generic_type of TCM_READ_WAIT : constant is 1;
    attribute mti_svvh_generic_type of TCM_WRITE_WAIT : constant is 1;
    attribute mti_svvh_generic_type of TCM_SETUP_WAIT : constant is 1;
    attribute mti_svvh_generic_type of TCM_DATA_HOLD : constant is 1;
    attribute mti_svvh_generic_type of TCM_TURNAROUND_TIME : constant is 1;
    attribute mti_svvh_generic_type of TCM_TIMING_UNITS : constant is 1;
    attribute mti_svvh_generic_type of TCM_READLATENCY : constant is 1;
    attribute mti_svvh_generic_type of TCM_SYMBOLS_PER_WORD : constant is 1;
    attribute mti_svvh_generic_type of USE_READDATA : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITEDATA : constant is 1;
    attribute mti_svvh_generic_type of USE_READ : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITE : constant is 1;
    attribute mti_svvh_generic_type of USE_BYTEENABLE : constant is 1;
    attribute mti_svvh_generic_type of USE_CHIPSELECT : constant is 1;
    attribute mti_svvh_generic_type of USE_LOCK : constant is 1;
    attribute mti_svvh_generic_type of USE_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of USE_WAITREQUEST : constant is 1;
    attribute mti_svvh_generic_type of USE_WRITEBYTEENABLE : constant is 1;
    attribute mti_svvh_generic_type of USE_OUTPUTENABLE : constant is 1;
    attribute mti_svvh_generic_type of USE_RESETREQUEST : constant is 1;
    attribute mti_svvh_generic_type of USE_IRQ : constant is 1;
    attribute mti_svvh_generic_type of USE_RESET_OUTPUT : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_READ : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_LOCK : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_WRITE : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_CHIPSELECT : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_BYTEENABLE : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_OUTPUTENABLE : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_WRITEBYTEENABLE : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_WAITREQUEST : constant is 1;
    attribute mti_svvh_generic_type of ACTIVE_LOW_BEGINTRANSFER : constant is 1;
    attribute mti_svvh_generic_type of CHIPSELECT_THROUGH_READLATENCY : constant is 1;
end system_0_cfi_flash_0;
