// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UFi/ONQXP5SVm68pPfyt96CDwaJYrhue/JxdXC55UE7lOH52ELwitP0qe5vdQkyu
T0XvgHYWcHbpWB3Ll7WptJL8R7/p+rU5EVUCq8W40hzw4hDR8VqdYW252jUaOAq3
NSWq1H/2JXeqiny9jp6H97VhSzkP+STHEdMr6OMqsLI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6096)
LyHdKkxL9Hsgi9CwwzB4sjWY9bP0TCqGUZdsxR9YNK1XqXMnfpZP/lA2DAi5FfFs
rUX61+iHrNduIX7wNtwhiHaDf/oc1MQIYGuXCNcwxAYphLvoxY2d/GmRziDTGV8t
tUCX2V95gfOw3DVfiZy0P/e3kF5I6GVAfRTx6RpSTD92qjOzXthF4ti0fHzMc44/
tG7zrJRXkIl3ofqH34F9/w0O3HeXbRUyqAPZkbfRDSLBZXQ6po9AbYRaqfRxqxGW
Yi5J3X7aj1nuinn1zGDwu/tHT/4C8Q603u6/vLiFclQnZj6KGCFuAQmu6MccbPSR
pEZsrqqtSWkol4yvaxsMHMzsshKiZeRoRnwyX2CQL6C0R+8bifM1n+mxFl+9Kg5t
5OQFdsbMx+TNeWytK0dOsFOBOJ1zNCri3KSi0XnuZenG4i/hLGzmIsbHIloGxNAo
pPx6QNQLS9iR/NoaOKtCurt7BSLIuESnFwOzggz/A+aHwGkYfQMoCW8WllGNKa/f
d1TI9RfQLF2lKQ3OwEwSMosPQA9w1yXRp8X8msMMzdqWB1qwgLWHvuPLKlRwVIQt
T2Whbjzp9zGr3C/NVictdoRGolLBNIXU2sIyADw/yqtJT3NTTlW3BsWeTLbn0Ynd
xD4bpJMD/yPltu/JdEUZDMODSQZROYgEf9HsetUca5z+cHZI0naDrD+h/uUsFIAv
WCad1/fR5Za25I6c5tOBEGg9HR9+hr2Gck38qiHBKC6nhQssqocGRh7raXZld9mS
gqRcHooS6CWpvSA49PFy0+RCqDDgMHAEqnhcZt/aWhyAJ0zfMVF/wG5KL9OxS9SZ
ZtfC9H5jZXvIfryFzs6j741woLuR6JRd/GV0jVbe91Lvm3popSVQkRgHYi03rmdf
/9FPOMVF5VNcurmk6r3ITNjiuRbO5ha5G21yFfIsb5C25O68CV1YPOgaQ/i4Ssj0
CkcagZJHh2p4oKhJtFdI29TKOaxSgtavKnx58hqDkRQlgFcNTHBylOa79zjT4+Hv
nI2wsjV1d7tmaM9op3pNK4ReQq+T25Vpod9tysUhos51QkgtVWXYGHP+O7ZngCZT
OyNWbZrwOxgJpdI8TVnnmElJNJwlzm/myDlE8vnJ/LRspGvcO2Ht2y0RzPLpcm01
xfLhTKzkzd0x7mUXF368GAoI7iICrLXm5lYDImMbbY0YJ2H5mJSrURaHywNc8gi1
5v0JVRHBi+MHhdW4Z5eAnIvsyePeoveHn//5ZimWPwNM0Ey2dsZICysoyYSI4mJ3
rRGkWtwOY/MubibCQdsIpeBcN0ArZ2pgsIet6zL7OwRN72wjDegFNRmWu7JeCv0k
kICohuuybUxR7WfQQAhijCwj1bwTE7mazcuiTmKjsPFn4u8KNqnhOL6u7KLOT8Km
rbDnCZk37jdSTIQohRmSIIXVGJ6WvnRS/AHo6ECg6+JERKDyhQ9lLlz82PJXjjzQ
TzmUMVHAqD4tkdVlMkLQxuCtRBbB5J1jtwRIb2qwexrwklEOJzFxNZkEB1FBkcf3
AVUfu5p/Wf43SjKJq4TFWqaQa0k6uEjoPAYSO8jLW/6kQbOCDBMxc+FReNp1i+18
WLYQL8fGbyqhgOuiCLyx4Pta3OfUc1Imw0Sz5HGlUsz5rmAjKcZrwEZKTN3YNWil
dkFLoGJYIBlsyXjCZoStTJ87tw8D+rPi7A5UpCGRyxRnwYeCIceE8CG1/Dh9wqsK
9lKijGpFmzjXNMUY2eWJ6xDmEa8+0SMql8ZVYP+716BeRmXlPDDtqOCJqY3LLOE6
MCu8eAG7uLYkvHQFLDdncE7n+B8sNzK+lXEnhFNG1f0k2/6Oa7sqt7H+4lsnaUSc
egVykLBJBvrDX3byGnCBdnMukkT+F/Qwa01DsC9ktUEDM+K4Zo1Kb5SrE7CEuubO
axQg99R5q/kgxC81Fkd45Y4GTaHFHlTLDBIuCeQGDDzikRQ7wRa3xC5/RbABCJwq
mLBUmxiUDvNzixNDRR/2A8fbXwEoL6mtjyCNqfTPw+oD+o4AbNpv98ov2z2wU9we
PVMr2fEA3FuIGPlEBB0H1t8VFmo7QQuRu8xN1tGlxyAooKoIK/kR3Ri2EpUUwVE/
NgNPJj5DRUFW++UPAaXVDAWjo7DGVmP5mxnNCIxFUzkytw53zncXtJgZImjH8rFH
mkTK+BAQpeN2HGEQfeUJ3i2xrogku832CS3V9x9C0WYqSDmaF1/B50mTgoHq54Oq
FYrQ68jsSVFNrhQcz9ODf6z8LwE/txdrTvGWBqxBZ4ODcHzU2diTRjr2MKhvYbw2
YnhPz63834aWFEb8r2ZNeV4MyEIbB3wBd4GplP+vXEcNd+a352bRBeN+XbybKGdS
TZ0bDOkG+0yDtK0eZQmZegAL3MCu3JKSc+w1znmE4GVkgY1ITy8fI3mgR2KP1cp5
BtO42Tv364bT41a+oVZc3Axv199/ORBCZlUJbzxScpIhiOXUcS0B4V1URDPbXe8J
6hvuWaAEcftcpuQWgteyFZWev+M97pv2KN/E80b82EVnACbiQkzRivM0jD4nXske
KAS9uZLij1I1UNGHrLHqkKg89NjT0NYEx3whHj1dL0z6EON7Wp8s4T8Xt9Ly2mF+
BWdGpuz4P66hfPNqoIt87fesHylkiMgGTmoV6RL9DNT9ifvaairzEvGnzaXRsihu
RaYMHr4aTe3DBOajI6sf8EAbnP+pbcKGfSB8URcX5RzCIzQGhnYa2YYzP2QqCiFf
wu6zcGUiJGhRXV57GA/ZFW88GoL0ECoue1HV/wxpCke5FZXdiMeIoV9/76Kt4dAp
o7XeUDhQr04gjVK7c1iLO0xsATSevqTyuXApPWSZBS2D3enMk+CmHDHSbNPbO9dx
g8cavFfAzR8g3eOfaRqoxvrwxc7mbZy6tFHTXfwBnlfOKQ3Dn2Sg/FBDV4FySa1r
iuKpSqLwGtjtBwNBhJygDo2kltqqx/77cZaOjbwaXRY8pPCZ5RZB1RppuoeDZ4NU
2lWbcZExJXNG390N0i+LC0KCz3n7iMTNpjA21T0GtlvquwJEMBJJ8Z9i30gvqw6d
dgD1UqPapyWEp/fS+lkquJbpcHgTRGQeOr2gLSXLX5IQz2gbINoZY70YWoE2K2TZ
NpL9Qcl/XX5RzVCYiskXwBmK0RobOWeUs3Ho5QCTHYLiQNrYZE1DNO6vhT5fJ3pZ
2hjQO9coTP37CJqvHCem0pQv5x+FR4Aw5VmuOGNl1JAxHh2TX/74WsLWP36lNOSt
njHNg3SnlRR8EQ3hrUu22EE6ZQdWNH8KzIMxTfzBsB3Y1q4uAXFe6N4fBNn+IMy3
wOgUJHq2s44megFiwXGs5q2+UK9APJEIz3h764rLphSQtGjxq4/t6zredXZnJnG8
BL13edAVFIXvJI78ATE8l3myK5qLhh7ZMOXoji+HTnLMPzZQc0DAr4+4VbesP0X1
Jr4n7zwdFwhn4YrrTnq0L5ZZoPXQN/Lg3tcGcK5nYCUCs9l7A/75yGSSwdP5YRRy
RbPXYvpt4Q9yVeneZfxQB2vOqaSrqLrI+4rNmXATVW+SOPuzdVG0YlpLkOPTN2KC
eDD9k+3dVR8SDX8ABFTan3M5KhtJr/uTRh3oel3mhhNjyY+TNxfZ/j3lxylRi2ja
AY2XKGKsx80K9UvOcitpOwnUdmrh7asFePF/pdj0dcDvdE1vFFQEpsKBrS37kv+J
SqRSIKJjq3p+PZU3prSVm56KjHOVkSAhcyKD5gGXdkevSgsP68S+yP36Lcv56dcS
N69coXq255x2xoXRQ1MCGOFvFCnvG9iX3FbcBK91ZjcMjab9HYmqltIbwP1TXtoF
UYIlVfXKZdQ7M/UsU/gwErhZ5uftCg/qJdm+GatKdPtzzcNEWwrNWPoKaf7CfPoh
1/T0pv8tiW25UvJnWkPAB8rMIUsg1qFXrJr65vAdZm/K5sobM2++41VuEwDF4JZx
oWHW95u7mz+oV1y0mXLJ51C5XJysF8etpNSDl1DQn2cSGhrUjN2mb8dxQH2gL6Sg
VrOQlBQiFa5jfCwUrtIKDNSTTNKgUnjLPftQjsvCtSoj7KjS42OI5IpHnGcAve89
wuks70DXkGq8JKkqPqSzW4m6QMiH7L27sB/fc3aWdD3xZBsK4Xw5l3UhSqM7sdxh
rAl1gzsPehRr1gwMcv7MQFYrSY0KFUNlWkb+6OiMViR4SAVVZWV6Mw4QvfUsSB3b
5UZV7FzhQjTZnJeMTlKNrKJgfCt1M7j77Bsb5FdJLjqPi1TzVIiyK8FJkIVsGOzO
W1oaeIpYSm46oSynpU/DjTp2gUs8RR/82PKCWS5VasYhJCfZYX2AjGLYylJR0Gnr
w5QsrTDkUajJpbp28BwbXmN9/R63bV6mkaEOIx9g6X1lfOLRbi1jcAecJu9/3iCk
CllRPy6sFfSAZWZXrORwwpS5Tu2zwgqs/ktyCeUDeRPBbxAf1LXgpAjsWC3+V1jH
8HB6T5BWGyRJSJcn7TjIVgd5g6mLfkhZLcQ4PTIfCdJZoiOwt9k0UA/dsgpYQaI+
u0YlRPm+ILFQxn/jfsCNABHVy2VYjG+NdTIgD8zRXm/0psVM5pg+LUT2b9w3wLv3
PAwqktT60IFD/CIKzzvwfyzMesXmjPUSRf90vT0dVa+cey8BcJtn3Bu/wlMcUnYs
yszVEHxTTFTbQh8z7ccAI6hWK6SEhVCa/oOyIjK4/HDSuQBFhjX/rnwnchYEE+Uf
Ul+2nMexzgcemXfHcB0euX1TA5QnpKApIhNoCEeCrwBfdgqwFcMusI9whCbBdExO
ELGs+xJXdSmwChH9jF0hytZcEEJ7ddct0cEqUXpk+h7RrsG/tUTuRuO2XPHXBIld
wEgX2fJJzV4C/dg/5/oMv7JMke+pZaohUyd1C2sWfHm7gx3HbX4a6dH7QwJiuwHf
AiSRPXUCDzZugMiY4vW9VM+69TJk5/TraAw48LBsgvQEgIbpMe1ZeCIbbdh1buqX
huQiGuzFhRB6HRJ+8qu5epfpt1mvQyW2hgpKwy3x6URsPkikSgKqF+nXTJtY4Pti
honssJswCqzQhqH9IkWVHSJWNlCWV15LZ4I/Z/Xa+H76dwZ1p/1O0BA2/DuMHz81
NUgs6P/IxL0PIYMFL/G87x9vzqxQF5ux4k5P/fTZp3J/kLYZmHG0Wv7YyoWD1IZI
Pqm9GkHUhKA9XFDi2At1rQOGEESKQmbshuohxqjBGu3ewfFJQ4a9aN1gpyhNNeZf
pRhMUbdhn/bin7qMHjhFKmaUM7QxwsjYhqEI/GsTzwOTyyUARJ0Quuh3gU2VPiO/
6KgjmbvoShZ23a+5znN6TkjrH+y+rMUixwtEZxAO+Y2BxoPyTdG4SHM72Y6c54GY
FiixF1UCeeygD+ZdnVlznvLSsOyIFtWpJz+CtA1E/PW6Kp/rON0dlm63cbZVzMYu
9fl+MMs9t8HJJH+B6SnfoKcPILAFbInZir/unKHPcP8nEgrItfqD3hl0/Pq5+oJm
6C0MVienMFvNARuvtppJg4Yghp9hY0rQB8/BOV36Yu8qC0o1FKy8+ODoz44tguC9
/QFT9k2lbeKJleeOk6jXlLngOOWROICchVrHI3qKXT6CTz4MJ9QNf2E5zW8dWY71
iXfUl3wFO0D7czisIHCuqIbjKR3dnbTmABAErHudOE5Zt52atPS9KbDW62aCqZ/L
SeC89q3o6Hr2AiYrc308EbxyHU2r9Ijjo1zFZ18UaxBkDPBef+amEbObyIORf76N
qTPc1C4L1Yd0q4ynjJFQF062KdAWCE9NVdm+3H8E5BoySZ4JS6GYNO7/y2EAvimB
PElo0K7KZTsO4P1M+NnH/8j7Du6s9q+9XWGakKNYaeuC5SSJurewxyhYjucGSFMg
8lMkbx3g+xMvwIiG/S7tPujrFw45tXLFwrs6Da44ZJ11DbUaORTNw7nbUriiACc+
2DMQh6IMlDiwrvpIhb6qhoZ/HC0ckIWbWY4XFIuoSlmzt0fk9BRj6K/YtjHbK2nH
j9XLMq+lnZQ/ldeWKE9MLK+GcZ4Iei7J1GpIA3ZK2qdujPNRTGZddHHLt2aUYKza
vdjMXliKSFexqoPgOGQMhxuT0eQOY3jLmrb8MlDXsFzVgUEiE7QDMAthy/9Y0Jp4
59njZYHWYlM/EFwHZOhd89YfIJBZhjCJH4Hxb+OTeqvE0aQzmhrtMHAS7u03DMsq
M63PaSIyKB6SuLN3eOZIPIOXwtkOfIOdhVLlk/wa9iEPjyEGT0clUIKMJ4fHGyHN
B64vAzX+WwfL63DMeOGKP2zQmuoVqNfhesNDn1avzRAa7iox+L/yjgW8IjLIwU9V
3AjGTwkHUZkG6o71BFxOhl4sQ9bt9JonqUs5p0kDi+MgCOoMAniASfyNJjO1kF5E
TS0zHlM2rvyzMuxTLtlUqFs0VVlya/3qgFZMD0/iezdQ9S6Hnk7cBBv5zXC48LbM
PE349wuOA+GUeMB2XHAAu1s2DZfYIESWQPVT5AHMpo8eWEaegTxSlx5t5nffgymU
ZpGrHv7E5qG3fUdSKQ6E+KZzxGPYl9x3ISHYGCNCf4FhXnZbu8Ek3d7a9z92r0hT
QbwASaHJnAZZsnJjJTpPhIvXeW2Vgs8EmjpXa5LHNfy1dzZbvdfKrs+4Yb/WFo0k
Fk/uSoIhtG4TuuYfJWCEtouCzaFeF2wgJVf110nbNL2RETWzBdhqTfuvYAn8PPa1
IPOAZCD7G9am/bXqMs9OK/oU9N0Ee5lfjL4Ywl3y6y/DyMCgGEGmUpqoYLybR9Jy
pNHPQBvYL01UPWe2ryCIiIY08EEXvn2XryU/pr899jP0hkBKp/pHVehFbY25BjzB
sb+AwvrT1cIMO/AytHujuE9H4GJMOR3UVKxVyMouotGqh/s8pFbNni9tnY4uCiH/
0+q+waPbE4zXXHr+8JRAkFXkIbYzGDblGhF8sOanERN2sQbwTQmi0wskf7Mi2P5w
tfPTB87YBH55O1wM67GqyahEvp5pqPSNcglAnNt12WY3zFkpHuHojnk8c0KxdzrY
VwNPXnKrqBx2KS+0B8BZgywKo27xYszkvPWT4UVGQ75Pl5R+A05YkkpOQM6gn287
LLI5UQndRgZdENi/AxZAUczcQk6P++k0aQSkm/E+N1BVwJdfx+niX52XezwZA0wC
ImVughFMydTp33tSAMWFszhh/Qqwoee9OBMn0uUPK5fHY6bEHDZlnAWDCspEUMdN
O0ZvvBH6ZJpfjsjamo9J5yll9wYsMAdFyvJsL4yCEx4/+nJIDBr427op7or8fwaG
8HIGt06QzQgrCFyaxjjIWiflC1ZLESgjxqZhBDM66OriKUbqlhfnqLp4gw73GXF9
45V6nS9MSZ3AM0DwbWUmE9t+CZmk3vc09T9xreqGy/W175rds1IsYfMkf0CNlX2b
nVPF6Gt2MWhSBCSOGCaK+qBwzwJYdyoZX01H9KVNhOhMRAyivX9wRBWp9VURz7MJ
oRraq4zbwY/zd0t2lJFp4DwALP2tJEI+X1ceZX88Jhbt6bq5DhC6qLkMC6Nr1umc
hc1DUKFvKLIpyyc66CLO19Rk4s+UVFQf/QeipEUtjfpUqZYLfw52/+vkkZxkbMhJ
kYnUjaHL2dcblmngmNpnAAOFyu77fkyHCo6pO3ECXS+v5DZfgrlBA+ixzHzx6WNw
ddEMKEOCkyHRuTIb+rwZ/1Kum5Mjc3rR6v5yBjiedaxyvOaMGFCfGo+nMfkJ4QXo
AGNppJ2FyKUFyOjMOyHzOXwWH8d2CHgkHgEP6LOVTbokajGSsDxjVlr0PFY3eXr+
CYKURtJ9wbyqzFJCqhX5AU7DrzluS/i0iyTBsyMtGI6bv8OyE4re76hXleGE6pyd
zaolMQAbHjTxZbdTlKvJYwMzVAkrBX5SSuYVJIGaZW+lJBF4PaUI12kllo3d+jdi
Rc4HHtscst5v/OXUEQL62svpV8eKEtd6Iz916NcRlgkahF1LEfqHxOzLOx4SKdYw
sjFqrFxyW4kp4zpqHExeOqc3/s16bsHAuVUK6kPKgGalaDYs4zVm5SS7e3dUiZ4U
yaeRdbNNg1dRZU6xIAELVyCLxMw4ht4ol23pGWHZnDRoPg6vFji4/tmnFDESBJu+
`pragma protect end_protected
